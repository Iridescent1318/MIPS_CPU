
module DataMemory(reset, clk, Address, Write_data, Read_data, MemRead, MemWrite);
	input reset, clk;
	input [31:0] Address, Write_data;
	input MemRead, MemWrite;
	output [31:0] Read_data;
	
	parameter RAM_SIZE = 256;
	parameter RAM_SIZE_BIT = 8;
	
	reg [31:0] RAM_data[RAM_SIZE - 1: 0];
	
	assign Read_data = MemRead? RAM_data[Address[RAM_SIZE_BIT + 1:2]]: 32'h00000000;
	
	integer i;
	
	initial begin
	    RAM_data[0] = 32'd306;
        RAM_data[1] = 32'd328;
        RAM_data[2] = 32'd738;
        RAM_data[3] = 32'd38;
        RAM_data[4] = 32'd901;
        RAM_data[5] = 32'd56;
        RAM_data[6] = 32'd301;
        RAM_data[7] = 32'd705;
        RAM_data[8] = 32'd293;
        RAM_data[9] = 32'd593;
        RAM_data[10] = 32'd923;
        RAM_data[11] = 32'd370;
        RAM_data[12] = 32'd477;
        RAM_data[13] = 32'd353;
        RAM_data[14] = 32'd781;
        RAM_data[15] = 32'd865;
        RAM_data[16] = 32'd979;
        RAM_data[17] = 32'd519;
        RAM_data[18] = 32'd952;
        RAM_data[19] = 32'd748;
        RAM_data[20] = 32'd501;
        RAM_data[21] = 32'd514;
        RAM_data[22] = 32'd690;
        RAM_data[23] = 32'd389;
        RAM_data[24] = 32'd68;
        RAM_data[25] = 32'd291;
        RAM_data[26] = 32'd343;
        RAM_data[27] = 32'd559;
        RAM_data[28] = 32'd501;
        RAM_data[29] = 32'd274;
        RAM_data[30] = 32'd862;
        RAM_data[31] = 32'd109;
        RAM_data[32] = 32'd457;
        RAM_data[33] = 32'd499;
        RAM_data[34] = 32'd381;
        RAM_data[35] = 32'd991;
        RAM_data[36] = 32'd242;
        RAM_data[37] = 32'd795;
        RAM_data[38] = 32'd711;
        RAM_data[39] = 32'd140;
        RAM_data[40] = 32'd993;
        RAM_data[41] = 32'd793;
        RAM_data[42] = 32'd525;
        RAM_data[43] = 32'd293;
        RAM_data[44] = 32'd280;
        RAM_data[45] = 32'd84;
        RAM_data[46] = 32'd32;
        RAM_data[47] = 32'd667;
        RAM_data[48] = 32'd672;
        RAM_data[49] = 32'd462;
        RAM_data[50] = 32'd109;
        RAM_data[51] = 32'd972;
        RAM_data[52] = 32'd984;
        RAM_data[53] = 32'd435;
        RAM_data[54] = 32'd484;
        RAM_data[55] = 32'd986;
        RAM_data[56] = 32'd404;
        RAM_data[57] = 32'd531;
        RAM_data[58] = 32'd386;
        RAM_data[59] = 32'd302;
        RAM_data[60] = 32'd521;
        RAM_data[61] = 32'd411;
        RAM_data[62] = 32'd94;
        RAM_data[63] = 32'd346;
        RAM_data[64] = 32'd232;
        RAM_data[65] = 32'd78;
        RAM_data[66] = 32'd771;
        RAM_data[67] = 32'd929;
        RAM_data[68] = 32'd332;
        RAM_data[69] = 32'd588;
        RAM_data[70] = 32'd781;
        RAM_data[71] = 32'd687;
        RAM_data[72] = 32'd982;
        RAM_data[73] = 32'd436;
        RAM_data[74] = 32'd269;
        RAM_data[75] = 32'd804;
        RAM_data[76] = 32'd806;
        RAM_data[77] = 32'd829;
        RAM_data[78] = 32'd16;
        RAM_data[79] = 32'd516;
        RAM_data[80] = 32'd747;
        RAM_data[81] = 32'd454;
        RAM_data[82] = 32'd3;
        RAM_data[83] = 32'd321;
        RAM_data[84] = 32'd473;
        RAM_data[85] = 32'd190;
        RAM_data[86] = 32'd924;
        RAM_data[87] = 32'd511;
        RAM_data[88] = 32'd652;
        RAM_data[89] = 32'd49;
        RAM_data[90] = 32'd966;
        RAM_data[91] = 32'd802;
        RAM_data[92] = 32'd492;
        RAM_data[93] = 32'd977;
        RAM_data[94] = 32'd81;
        RAM_data[95] = 32'd364;
        RAM_data[96] = 32'd953;
        RAM_data[97] = 32'd564;
        RAM_data[98] = 32'd980;
        RAM_data[99] = 32'd169;
	    for(i = 100; i < RAM_SIZE; i = i + 1) RAM_data[i] <= 32'h00000000;
	end   
	
	always @(posedge reset or posedge clk)
		if (reset) begin
		    RAM_data[0] = 32'd306;
            RAM_data[1] = 32'd328;
            RAM_data[2] = 32'd738;
            RAM_data[3] = 32'd38;
            RAM_data[4] = 32'd901;
            RAM_data[5] = 32'd56;
            RAM_data[6] = 32'd301;
            RAM_data[7] = 32'd705;
            RAM_data[8] = 32'd293;
            RAM_data[9] = 32'd593;
            RAM_data[10] = 32'd923;
            RAM_data[11] = 32'd370;
            RAM_data[12] = 32'd477;
            RAM_data[13] = 32'd353;
            RAM_data[14] = 32'd781;
            RAM_data[15] = 32'd865;
            RAM_data[16] = 32'd979;
            RAM_data[17] = 32'd519;
            RAM_data[18] = 32'd952;
            RAM_data[19] = 32'd748;
            RAM_data[20] = 32'd501;
            RAM_data[21] = 32'd514;
            RAM_data[22] = 32'd690;
            RAM_data[23] = 32'd389;
            RAM_data[24] = 32'd68;
            RAM_data[25] = 32'd291;
            RAM_data[26] = 32'd343;
            RAM_data[27] = 32'd559;
            RAM_data[28] = 32'd501;
            RAM_data[29] = 32'd274;
            RAM_data[30] = 32'd862;
            RAM_data[31] = 32'd109;
            RAM_data[32] = 32'd457;
            RAM_data[33] = 32'd499;
            RAM_data[34] = 32'd381;
            RAM_data[35] = 32'd991;
            RAM_data[36] = 32'd242;
            RAM_data[37] = 32'd795;
            RAM_data[38] = 32'd711;
            RAM_data[39] = 32'd140;
            RAM_data[40] = 32'd993;
            RAM_data[41] = 32'd793;
            RAM_data[42] = 32'd525;
            RAM_data[43] = 32'd293;
            RAM_data[44] = 32'd280;
            RAM_data[45] = 32'd84;
            RAM_data[46] = 32'd32;
            RAM_data[47] = 32'd667;
            RAM_data[48] = 32'd672;
            RAM_data[49] = 32'd462;
            RAM_data[50] = 32'd109;
            RAM_data[51] = 32'd972;
            RAM_data[52] = 32'd984;
            RAM_data[53] = 32'd435;
            RAM_data[54] = 32'd484;
            RAM_data[55] = 32'd986;
            RAM_data[56] = 32'd404;
            RAM_data[57] = 32'd531;
            RAM_data[58] = 32'd386;
            RAM_data[59] = 32'd302;
            RAM_data[60] = 32'd521;
            RAM_data[61] = 32'd411;
            RAM_data[62] = 32'd94;
            RAM_data[63] = 32'd346;
            RAM_data[64] = 32'd232;
            RAM_data[65] = 32'd78;
            RAM_data[66] = 32'd771;
            RAM_data[67] = 32'd929;
            RAM_data[68] = 32'd332;
            RAM_data[69] = 32'd588;
            RAM_data[70] = 32'd781;
            RAM_data[71] = 32'd687;
            RAM_data[72] = 32'd982;
            RAM_data[73] = 32'd436;
            RAM_data[74] = 32'd269;
            RAM_data[75] = 32'd804;
            RAM_data[76] = 32'd806;
            RAM_data[77] = 32'd829;
            RAM_data[78] = 32'd16;
            RAM_data[79] = 32'd516;
            RAM_data[80] = 32'd747;
            RAM_data[81] = 32'd454;
            RAM_data[82] = 32'd3;
            RAM_data[83] = 32'd321;
            RAM_data[84] = 32'd473;
            RAM_data[85] = 32'd190;
            RAM_data[86] = 32'd924;
            RAM_data[87] = 32'd511;
            RAM_data[88] = 32'd652;
            RAM_data[89] = 32'd49;
            RAM_data[90] = 32'd966;
            RAM_data[91] = 32'd802;
            RAM_data[92] = 32'd492;
            RAM_data[93] = 32'd977;
            RAM_data[94] = 32'd81;
            RAM_data[95] = 32'd364;
            RAM_data[96] = 32'd953;
            RAM_data[97] = 32'd564;
            RAM_data[98] = 32'd980;
            RAM_data[99] = 32'd169;
			for (i = 100; i < RAM_SIZE; i = i + 1)
				RAM_data[i] <= 32'h00000000;
		end
		else if (MemWrite)
			RAM_data[Address[RAM_SIZE_BIT + 1:2]] <= Write_data;
			
endmodule
